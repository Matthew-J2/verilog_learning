module mod_a (input in1, input in2, output out);
    mod_b inst(a,b,out);
endmodule
