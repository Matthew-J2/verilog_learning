module hello_verilog_2 (
    output zero
);

  assign zero = 1'b0;

endmodule

